library ieee;
use ieee.std_logic_1164.all;

ENTITY REG_7 IS
	PORT(
		DIN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		CLK : IN STD_LOGIC;
		DOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END REG_7;

ARCHITECTURE BEHAV OF REG_7 IS
	BEGIN
		PROCESS (CLK)
		BEGIN
			 IF RISING_EDGE(CLK) THEN
						DOUT <= DIN;
			 END IF;
		END PROCESS;
END BEHAV;
