LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

package types_pkg IS
	CONSTANT N_PARTIAL_PRODUCT : integer := 17;
	CONSTANT PARALLELISM 	:	INTEGER := 32;
	
	CONSTANT STRT_COL_L7		:	INTEGER := 24;
	CONSTANT NUM_HA_FA_L7	:	INTEGER := 18;	--there are 19 adders, so from 0 to 18
	CONSTANT END_COL_L7		:	INTEGER := 42;
	CONSTANT NUM_OP_L7		:	INTEGER := 16; --there are 17 operands, so from 0 to 16	
	CONSTANT DEPTH_L7			:	INTEGER := 3;	--there are 4 HA and FA layers, so from 0 to 3 
	
	CONSTANT STRT_COL_L6		:	INTEGER := 16;
	CONSTANT NUM_HA_FA_L6	:	INTEGER := 34;
	CONSTANT END_COL_L6		:	INTEGER := 50;
	CONSTANT NUM_OP_L6		:	INTEGER := 12;
	CONSTANT DEPTH_L6			:	INTEGER := 3;
	
	CONSTANT STRT_COL_L5		:	INTEGER := 10;
	CONSTANT NUM_HA_FA_L5	:	INTEGER := 46;
	CONSTANT END_COL_L5		:	INTEGER := 56;
	CONSTANT NUM_OP_L5		:	INTEGER := 8;
	CONSTANT DEPTH_L5			:	INTEGER := 2;
	
	CONSTANT STRT_COL_L4		:	INTEGER := 6;
	CONSTANT NUM_HA_FA_L4	:	INTEGER := 54;
	CONSTANT END_COL_L4		:	INTEGER := 60;
	CONSTANT NUM_OP_L4		:	INTEGER := 5;
	CONSTANT DEPTH_L4			:	INTEGER := 1;
	
	CONSTANT STRT_COL_L3		:	INTEGER := 4;
	CONSTANT NUM_HA_FA_L3	:	INTEGER := 58;
	CONSTANT END_COL_L3		:	INTEGER := 62;
	CONSTANT NUM_OP_L3		:	INTEGER := 3;
	CONSTANT DEPTH_L3			:	INTEGER := 0; 
	
	CONSTANT STRT_COL_L2		:	INTEGER := 2;
	CONSTANT NUM_HA_FA_L2	:	INTEGER := 61;
	CONSTANT END_COL_L2		:	INTEGER := 63;
	CONSTANT NUM_OP_L2		:	INTEGER := 2;
	CONSTANT DEPTH_L2			:	INTEGER := 0; 
	
	type PP IS array(0 TO N_PARTIAL_PRODUCT-1) of STD_LOGIC_VECTOR(PARALLELISM DOWNTO 0);
	type TABLE_L7 IS ARRAY(0 TO NUM_OP_L7) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type TABLE_L6 IS ARRAY(0 TO NUM_OP_L6) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type TABLE_L5 IS ARRAY(0 TO NUM_OP_L5) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type TABLE_L4 IS ARRAY(0 TO NUM_OP_L4) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type TABLE_L3 IS ARRAY(0 TO NUM_OP_L3) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type TABLE_L2 IS ARRAY(0 TO NUM_OP_L2) OF STD_LOGIC_VECTOR(63 DOWNTO 0);
	type S_C_L7 IS ARRAY(0 TO DEPTH_L7) OF STD_LOGIC_VECTOR(NUM_HA_FA_L7 DOWNTO 0);
	type S_C_L6 IS ARRAY(0 TO DEPTH_L6) OF STD_LOGIC_VECTOR(NUM_HA_FA_L6 DOWNTO 0);
	type S_C_L5 IS ARRAY(0 TO DEPTH_L5) OF STD_LOGIC_VECTOR(NUM_HA_FA_L5 DOWNTO 0);
	type S_C_L4 IS ARRAY(0 TO DEPTH_L4) OF STD_LOGIC_VECTOR(NUM_HA_FA_L4 DOWNTO 0);

end package types_pkg;

