library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types_pkg.all;

ENTITY UNFOLDED_FIR IS
		PORT(	D_IN_3K : IN SIGNED(Nb-1 DOWNTO 0);
				D_IN_3K_1 : IN SIGNED(Nb-1 DOWNTO 0);
				D_IN_3K_2 : IN SIGNED(Nb-1 DOWNTO 0);
				H0 : IN SIGNED(Nb-1 DOWNTO 0);
				H1 : IN SIGNED(Nb-1 DOWNTO 0);
				H2 : IN SIGNED(Nb-1 DOWNTO 0);
				H3 : IN SIGNED(Nb-1 DOWNTO 0);
				H4 : IN SIGNED(Nb-1 DOWNTO 0);
				H5 : IN SIGNED(Nb-1 DOWNTO 0);
				H6 : IN SIGNED(Nb-1 DOWNTO 0);
				H7 : IN SIGNED(Nb-1 DOWNTO 0);
				H8 : IN SIGNED(Nb-1 DOWNTO 0);
				H9 : IN SIGNED(Nb-1 DOWNTO 0);
				H10 : IN SIGNED(Nb-1 DOWNTO 0);
				V_IN : IN STD_LOGIC;
				RST_N : IN STD_LOGIC;
				CLK : IN STD_LOGIC;
				V_OUT : OUT STD_LOGIC;
				D_OUT_3K : OUT SIGNED(Nb-1 DOWNTO 0);
				D_OUT_3K_1 : OUT SIGNED(Nb-1 DOWNTO 0);
				D_OUT_3K_2 : OUT SIGNED(Nb-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEHAV OF UNFOLDED_FIR IS

--COMPONENTS DECLARATION

	COMPONENT REG_7 IS
		PORT( DIN : IN SIGNED(Nb-1 DOWNTO 0);
				CLK : IN STD_LOGIC;
				RST_N : IN STD_LOGIC;
				EN : IN STD_LOGIC;
				DOUT : OUT SIGNED(Nb-1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT REG_8 IS
		PORT( DIN : IN SIGNED(Nb DOWNTO 0);
				CLK : IN STD_LOGIC;
				RST_N : IN STD_LOGIC;
				EN : IN STD_LOGIC;
				DOUT : OUT SIGNED(Nb DOWNTO 0));
	END COMPONENT;
	
	COMPONENT FF IS
		PORT(
		D : IN STD_LOGIC;
		CLK : IN STD_LOGIC;
		RST_N : IN STD_LOGIC;
		EN : IN STD_LOGIC;
		Q : OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT FF_2 IS
		PORT(
		D : IN STD_LOGIC;
		CLK : IN STD_LOGIC;
		RST_N : IN STD_LOGIC;
		EN : IN STD_LOGIC;
		Q : OUT STD_LOGIC);
	END COMPONENT;
	
-- Signals declaration
	SIGNAL b : coeff_array;
	SIGNAL D_STAGE_3K : data_array; -- DATA IN AND OUT FROM REGISTERS STAGE 3K
	SIGNAL D_STAGE_3K_1 : data_array; -- DATA IN AND OUT FROM REGISTERS STAGE 3K+1
	SIGNAL D_STAGE_3K_2 : data_array_2; -- DATA IN AND OUT FROM REGISTERS STAGE 3K+22
	SIGNAL POTATO_FF: data_ff; -- DATA BETWEEN FFs
	SIGNAL OUT_MULT_3K : mult_out_array; -- DATA FOR OUT MULT STAGE 3K
	SIGNAL OUT_MULT_TRUNC_3K : mult_in; -- DATA FOR TRUNCATION STAGE 3K
	SIGNAL OUT_ADD_3K : add_in_from_mult;  -- DATA FOR OUT ADD STAGE 3K
	SIGNAL OUT_MULT_3K_1 : mult_out_array; -- DATA FOR OUT MULT STAGE 3K+1
	SIGNAL OUT_MULT_TRUNC_3K_1 : mult_in;  -- DATA FOR TRUNCATION STAGE 3K+1
	SIGNAL OUT_ADD_3K_1 : add_in_from_mult;  -- DATA FOR OUT ADD STAGE 3K+1
	SIGNAL OUT_MULT_3K_2 : mult_out_array;  -- DATA FOR OUT MULT STAGE 3K+2
	SIGNAL OUT_MULT_TRUNC_3K_2 : mult_in;  -- DATA FOR TRUNCATION STAGE 3K+2
	SIGNAL OUT_ADD_3K_2 : add_in_from_mult;  -- DATA FOR IN ADD STAGE 3K+2
	SIGNAL ADD_IN_3K : add_in_from_sum; -- DATA FOR IN ADD STAGE 3K
	SIGNAL ADD_IN_3K_1 : add_in_from_sum;  -- DATA FOR IN ADD STAGE 3K+1
	SIGNAL ADD_IN_3K_2 : add_in_from_sum;  -- DATA FOR IN ADD STAGE 3K+2

	BEGIN
	
-- WE USED AN ARRAY FOR COEFFICIENTS IN ORDER TO BETTER USE PARAMETRIZATION IN THE ENTITY

	b(0) <= H0;
	b(1) <= H1;
	b(2) <= H2;
	b(3) <= H3;
	b(4) <= H4;
	b(5) <= H5;
	b(6) <= H6;
	b(7) <= H7;
	b(8) <= H8;
	b(9) <= H9;
	b(10) <= H10;
	
-- FFs

		FFs: FOR I IN 0 TO Nt GENERATE
			  FIRST_ITER: IF I = 0 GENERATE  
				  FF_IN:   		FF PORT MAP (V_IN, CLK, RST_N, V_IN, POTATO_FF(I));
				           END GENERATE;
							  
				LAST_ITER: IF I=Nt GENERATE
				  FF_OUT: FF_2 PORT MAP (POTATO_FF(I-1), CLK, RST_N, V_IN, V_OUT);
							  END GENERATE;
				
				INTERMEDIUM_ITER: IF ((I /= 0) AND (I /= Nt)) GENERATE
								FF_INNER1:	FF PORT MAP (POTATO_FF(I-1), CLK, RST_N, V_IN, POTATO_FF(I));
										END GENERATE;
			  END GENERATE;
	
-- INPUT REGISTER STAGE 3K

	INPUT_REG_3K: REG_7 PORT MAP (DIN => D_IN_3K, CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K(0));
	
	REG_STAGE_3K : FOR I IN 1 TO NT+1 GENERATE
					INT_REG: REG_7 PORT MAP (DIN => D_STAGE_3K(I-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K(I));
					END GENERATE;
	OUTPUT_REG_3K: REG_7 PORT MAP (DIN => OUT_ADD_3K(NT-2)(Nb-1 DOWNTO 0), CLK => CLK, EN => POTATO_FF(Nt-1), RST_N => RST_N, DOUT => D_OUT_3K);
					
--	MULTIPLICATIONS AND TRUNCATIONS STAGE 3K

		OUT_MULT_3K(0) <= D_STAGE_3K(0) * b(0);
		OUT_MULT_3K(1) <= D_STAGE_3K_2(1) * b(1);
		OUT_MULT_3K(2) <= D_STAGE_3K_1(2) * b(2);
		OUT_MULT_3K(3) <= D_STAGE_3K(3) * b(3);
		OUT_MULT_3K(4) <= D_STAGE_3K_2(5) * b(4);
		OUT_MULT_3K(5) <= D_STAGE_3K_1(6) * b(5);
		OUT_MULT_3K(6) <= D_STAGE_3K(7) * b(6);
		OUT_MULT_3K(7) <= D_STAGE_3K_2(9) * b(7);
		OUT_MULT_3K(8) <= D_STAGE_3K_1(10) * b(8);
		OUT_MULT_3K(9) <= D_STAGE_3K(11) * b(9);
		OUT_MULT_3K(10) <= D_STAGE_3K_2(13) * b(10);
		
		FIR_MULT_3K: FOR I IN 0 TO Nt-1 GENERATE
							REGS: REG_8 PORT MAP (DIN => OUT_MULT_3K(I)(2*Nb-1 DOWNTO Nb-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => OUT_MULT_TRUNC_3K(I));
						END GENERATE;
						
-- SUMS STAGE 3K

		OUT_ADD_3K(0) <= OUT_MULT_TRUNC_3K(0) + OUT_MULT_TRUNC_3K(1);
		REGS_3K: REG_8 PORT MAP (DIN => OUT_ADD_3K(0), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K(0)); --Da vedere

		
		FIR_SUM_3K: FOR I IN 1 TO NT-2 GENERATE
					OUT_ADD_3K(I) <= OUT_MULT_TRUNC_3K(I+1) + ADD_IN_3K(I-1);
					REGS: REG_8 PORT MAP (DIN => OUT_ADD_3K(I), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K(I)); --Da vedere
					END GENERATE;
	
-- INPUT REGISTER STAGE 3K+1

	INPUT_REG_3K_1: REG_7 PORT MAP (DIN => D_IN_3K_1, CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K_1(0));
	
	REG_STAGE_3K_1 : FOR I IN 1 TO NT+1 GENERATE
					INT_REG: REG_7 PORT MAP (DIN => D_STAGE_3K_1(I-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K_1(I));
					END GENERATE;
	OUTPUT_REG_3K_1: REG_7 PORT MAP (DIN => OUT_ADD_3K_1(NT-2)(Nb-1 DOWNTO 0), CLK => CLK, EN => POTATO_FF(Nt-1), RST_N => RST_N, DOUT => D_OUT_3K_1);
	
--	MULTIPLICATIONS AND TRUNCATIONS STAGE 3K+1

		OUT_MULT_3K_1(0) <= D_STAGE_3K_1(0) * b(0);
		OUT_MULT_3K_1(1) <= D_STAGE_3K(0) * b(1);
		OUT_MULT_3K_1(2) <= D_STAGE_3K_2(2) * b(2);
		OUT_MULT_3K_1(3) <= D_STAGE_3K_1(3) * b(3);
		OUT_MULT_3K_1(4) <= D_STAGE_3K(4) * b(4);
		OUT_MULT_3K_1(5) <= D_STAGE_3K_2(6) * b(5);
		OUT_MULT_3K_1(6) <= D_STAGE_3K_1(7) * b(6);
		OUT_MULT_3K_1(7) <= D_STAGE_3K(8) * b(7);
		OUT_MULT_3K_1(8) <= D_STAGE_3K_2(10) * b(8);
		OUT_MULT_3K_1(9) <= D_STAGE_3K_1(11) * b(9);
		OUT_MULT_3K_1(10) <= D_STAGE_3K(12) * b(10);
		
		FIR_MULT_3K_1: FOR I IN 0 TO Nt-1 GENERATE
							REGS: REG_8 PORT MAP (DIN => OUT_MULT_3K_1(I)(2*Nb-1 DOWNTO Nb-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => OUT_MULT_TRUNC_3K_1(I));
						END GENERATE;
					 
-- SUMS STAGE 3K+1

		OUT_ADD_3K_1(0) <= OUT_MULT_TRUNC_3K_1(0) + OUT_MULT_TRUNC_3K_1(1);
		REGS_3K_1: REG_8 PORT MAP (DIN => OUT_ADD_3K_1(0), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K_1(0)); --Da vedere
		
		FIR_SUM_3K_1: FOR I IN 1 TO NT-2 GENERATE
					OUT_ADD_3K_1(I) <= OUT_MULT_TRUNC_3K_1(I+1) + ADD_IN_3K_1(I-1);
					REGS: REG_8 PORT MAP (DIN => OUT_ADD_3K_1(I), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K_1(I)); --Da vedere
					END GENERATE;

-- INPUT REGISTER STAGE 3K+2

	INPUT_REG_3K_2: REG_7 PORT MAP (DIN => D_IN_3K_2, CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K_2(0));
	
	REG_STAGE_3K_2 : FOR I IN 1 TO NT+2 GENERATE
					INT_REG: REG_7 PORT MAP (DIN => D_STAGE_3K_2(I-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => D_STAGE_3K_2(I));
					END GENERATE;
	OUTPUT_REG_3K_2: REG_7 PORT MAP (DIN => OUT_ADD_3K_2(NT-2)(Nb-1 DOWNTO 0), CLK => CLK, EN => POTATO_FF(Nt-1), RST_N => RST_N, DOUT => D_OUT_3K_2);
	
--	MULTIPLICATIONS AND TRUNCATIONS STAGE 3K+2

		OUT_MULT_3K_2(0) <= D_STAGE_3K_2(0) * b(0);
		OUT_MULT_3K_2(1) <= D_STAGE_3K_1(0) * b(1);
		OUT_MULT_3K_2(2) <= D_STAGE_3K(1) * b(2);
		OUT_MULT_3K_2(3) <= D_STAGE_3K_2(3) * b(3);
		OUT_MULT_3K_2(4) <= D_STAGE_3K_1(4) * b(4);
		OUT_MULT_3K_2(5) <= D_STAGE_3K(5) * b(5);
		OUT_MULT_3K_2(6) <= D_STAGE_3K_2(7) * b(6);
		OUT_MULT_3K_2(7) <= D_STAGE_3K_1(8) * b(7);
		OUT_MULT_3K_2(8) <= D_STAGE_3K(9) * b(8);
		OUT_MULT_3K_2(9) <= D_STAGE_3K_2(11) * b(9);
		OUT_MULT_3K_2(10) <= D_STAGE_3K_1(12) * b(10);
		
		FIR_MULT_3K_2: FOR I IN 0 TO Nt-1 GENERATE
							REGS: REG_8 PORT MAP (DIN => OUT_MULT_3K_2(I)(2*Nb-1 DOWNTO Nb-1), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => OUT_MULT_TRUNC_3K_2(I));
						END GENERATE;
					 
-- SUMS STAGE 3K+2

		OUT_ADD_3K_2(0) <= OUT_MULT_TRUNC_3K_2(0) + OUT_MULT_TRUNC_3K_2(1);
		REGS_3K_2: REG_8 PORT MAP (DIN => OUT_ADD_3K_2(0), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K_2(0));
		
		FIR_SUM_3K_2: FOR I IN 1 TO NT-2 GENERATE
					OUT_ADD_3K_2(I) <= OUT_MULT_TRUNC_3K_2(I+1) + ADD_IN_3K_2(I-1);
					REGS: REG_8 PORT MAP (DIN => OUT_ADD_3K_2(I), CLK => CLK, EN => V_IN, RST_N => RST_N, DOUT => ADD_IN_3K_2(I));
					END GENERATE;
					
END ARCHITECTURE;
