Library ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

--SI POTREBBE METTERE NEI SEGNALI INSERITI DALLA CU UN QUALCOSA CHE SI PROPAGA LUNGO LA PIPE E CHE MI METTE LE NOP PER 3 CICLI (O 2?)

ENTITY Branch_Detection IS
	PORT(	ID_BRANCH_DET : IN STD_LOGIC;
			EX_BRANCH_DET : IN STD_LOGIC;
			PC_Write : OUT STD_LOGIC;
			IF_ID_Write : OUT STD_LOGIC;
			MUX_CU_BD : OUT STD_LOGIC
		 );
END ENTITY;

ARCHITECTURE BRAHVIOUR OF Branch_Detection IS
BEGIN

	PREDICTION : PROCESS (ID_BRANCH_DET, EX_BRANCH_DET)
	BEGIN
		IF ( ID_BRANCH_DET = '1' OR EX_BRANCH_DET = '1' ) THEN --HO UNA BEQ O UNA JAL CHE SI STA PROPAGANDO
			PC_Write <= '0';
			IF_ID_Write <= '0';
		ELSE
			PC_Write <= '1';
			IF_ID_Write <= '1';
		END IF;
		IF ( EX_BRANCH_DET = '1' ) THEN
			MUX_CU_BD <= '1';
		ELSE
			MUX_CU_BD <= '0';
		END IF;
	END PROCESS;
	
END ARCHITECTURE;
			