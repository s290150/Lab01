Library ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY RISCV_lite IS
	PORT(	instruction	:	IN		STD_LOGIC_VECTOR(31 DOWNTO 0);
			ReadData	:	IN		STD_LOGIC_VECTOR(31 DOWNTO 0);
			clock		:	IN		STD_LOGIC;
			reset		:	IN		STD_LOGIC;
			PC_address	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
			data_address:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
			WriteData	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
			MemWrite	:	OUT	STD_LOGIC;
			MemRead		:	OUT	STD_LOGIC
			);
	END ENTITY;

ARCHITECTURE structural OF RISCV_lite IS
--Component declaration
	COMPONENT sequencer IS
	PORT (JUMP_ADDR: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			PCSrc		: IN STD_LOGIC;
			PCWrite	: IN STD_LOGIC;
			clock		: IN STD_LOGIC;
			reset		: IN STD_LOGIC;
			I_ADDR	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT hazard_detection_unit IS
	PORT( RS1_ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			RS2_ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			EX_RD_ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			ID_EX_Mem_Read : IN STD_LOGIC;
			IF_ID_Write : OUT STD_LOGIC;
			PC_Write : OUT STD_LOGIC;
			MUX_CU_HD : OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT Branch_Detection IS
	PORT(	ID_BRANCH_DET : IN STD_LOGIC;
			EX_BRANCH_DET : IN STD_LOGIC;
			PC_Write : OUT STD_LOGIC;
			IF_ID_Write : OUT STD_LOGIC;
			MUX_CU_BD : OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT reg_file IS
	PORT(   RD_REG1	:	IN		STD_LOGIC_VECTOR(4 DOWNTO 0);
			RD_REG2	:	IN		STD_LOGIC_VECTOR(4 DOWNTO 0);
			WR_REG	:	IN		STD_LOGIC_VECTOR(4 DOWNTO 0);
			WR_DATA	:	IN		STD_LOGIC_VECTOR(31 DOWNTO 0);
			RegWrite	:	IN		STD_LOGIC;
			clock		:	IN		STD_LOGIC;
			reset		:	IN		STD_LOGIC;
			RD_DATA1	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
			RD_DATA2	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT immediate_generator IS
	PORT( 	immediate_in	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
			immediate_out	:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT execution_stage IS
	PORT( 	EX				: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			forwardA		: IN STD_LOGIC_VECTOR(1 DOWNTO 0);	
			forwardB		: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			PC_ADDR			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RD_DATA1		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RD_DATA2		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			IMMEDIATE		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			MEM_ALU_IMM		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			WB_WR_DATA		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			funct			: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			JMP_ADDR		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			Z_flag			: OUT STD_LOGIC;
			ALU_IMM			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT forwarding_unit IS
	PORT( EX_RS1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			EX_RS2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			MEM_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WB_RD  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			MEM_SW_BEQ : IN STD_LOGIC; --SE ABBIAMO UNA BEQ O SW NON ABBIAMO REGISTRI DI DESTINAZIONE
			WB_SW_BEQ : IN STD_LOGIC; --SE ABBIAMO UNA BEQ O SW NON ABBIAMO REGISTRI DI DESTINAZIONE
			FORWARD_A : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			FORWARD_B : OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT pipe_register_IF_ID IS
		PORT(	input	:	IN	STD_LOGIC_VECTOR(63 DOWNTO 0); --unconstrained array
				clock	:	IN	STD_LOGIC;
				reset	:	IN	STD_LOGIC;
				en_BD 		:   IN STD_LOGIC;
				en_HD 		:   IN STD_LOGIC;
				output	:	BUFFER	STD_LOGIC_VECTOR(63 DOWNTO 0)); --unconstrained array
	END COMPONENT;
	
	COMPONENT pipe_register_ID_EX IS
		PORT(	input	:	IN	STD_LOGIC_VECTOR(158 DOWNTO 0); --unconstrained array
				clock	:	IN	STD_LOGIC;
				reset	:	IN	STD_LOGIC;
				en 		:   IN STD_LOGIC;
				output	:	BUFFER	STD_LOGIC_VECTOR(158 DOWNTO 0)); --unconstrained array
	END COMPONENT;
	
	COMPONENT pipe_register_EX_MEM IS
		PORT(	input	:	IN	STD_LOGIC_VECTOR(107 DOWNTO 0); --unconstrained array
				clock	:	IN	STD_LOGIC;
				reset	:	IN	STD_LOGIC;
				en 		:   IN STD_LOGIC;
				output	:	BUFFER	STD_LOGIC_VECTOR(107 DOWNTO 0)); --unconstrained array
	END COMPONENT;
	
	COMPONENT pipe_register_MEM_WB IS
		PORT(	input	:	IN	STD_LOGIC_VECTOR(71 DOWNTO 0); --unconstrained array
				clock	:	IN	STD_LOGIC;
				reset	:	IN	STD_LOGIC;
				en 		:   IN STD_LOGIC;
				output	:	BUFFER	STD_LOGIC_VECTOR(71 DOWNTO 0)); --unconstrained array
	END COMPONENT;
	
	COMPONENT JAL_REG IS
		PORT(	input	:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0); --unconstrained array
				clock	:	IN	STD_LOGIC;
				reset	:	IN	STD_LOGIC;
				en 		:   IN STD_LOGIC;
				output	:	BUFFER	STD_LOGIC_VECTOR(31 DOWNTO 0)); --unconstrained array
	END COMPONENT;
	
	COMPONENT control_unit IS
	PORT(	OPCODE		:	IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			WB			:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
			M			:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
			EX			:	OUT	STD_LOGIC_VECTOR(5 DOWNTO 0));
	END COMPONENT;
	
--signals and types declaration

--IF STAGE

	--SEQUENCER SIGNALS
	SIGNAL JUMP_ADDR:	STD_LOGIC_VECTOR(31 DOWNTO 0); --PC + 4
	SIGNAL PCSrc		:	STD_LOGIC; --MUX SELECTOR BEFORE PC
	SIGNAL PCWrite	:	STD_LOGIC; --ENABLE PC
	SIGNAL I_ADDR	:	STD_LOGIC_VECTOR(31 DOWNTO 0); --OUTPUT PC
	
	--OR SIGNALS
	SIGNAL IF_ID_Write : STD_LOGIC;
	SIGNAL PC_Write : STD_LOGIC;
	
	--PIPE STAGE IF/ID IN & OUT
	SIGNAL IF_ID_input		:	STD_LOGIC_VECTOR(63 DOWNTO 0); --INPUT SIGNALS FOR PIPE STAGE
	SIGNAL IF_ID_output		: 	STD_LOGIC_VECTOR(63 DOWNTO 0); --OUTPUT SIGNALS TO PIPE STAGE
	SIGNAL ID_instruction	:	STD_LOGIC_VECTOR(31 DOWNTO 0); --OUTPUT OF INSTRUCTION MEMORY
	SIGNAL ID_I_ADDR 		: 	STD_LOGIC_VECTOR(31 DOWNTO 0); --SIGNAL USED AS INPUT IN THE NEXT PIPE STAGE
	
--DECODE STAGE
	
	--CU SIGNALS IN & OUT
	SIGNAL OPCODE	: STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL PREMUX_WB: STD_LOGIC_VECTOR(2 DOWNTO 0);	--forse sono meno per via della forwarding unit
	SIGNAL PREMUX_M	: STD_LOGIC_VECTOR(2 DOWNTO 0);--forse sono meno per via della forwarding unit
	SIGNAL PREMUX_EX: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL WB	 	: STD_LOGIC_VECTOR(2 DOWNTO 0);	--forse sono meno per via della forwarding unit
	SIGNAL M		: STD_LOGIC_VECTOR(2 DOWNTO 0);--forse sono meno per via della forwarding unit
	SIGNAL EX	 	: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL JAL_ctrl : STD_LOGIC;
	
	--SIGNAL FOR JAL_ADDR
	SIGNAL JAL_ADDR		: 	STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL WR_DATA_JAL	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ID_WR_DATA	:	STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL JAL_SEL		: STD_LOGIC;
	
	--REGISTER FILE SIGNALS IN
	SIGNAL RD_REG1	: STD_LOGIC_VECTOR(4 DOWNTO 0); --ADDRESS REG 1
	SIGNAL RD_REG2	: STD_LOGIC_VECTOR(4 DOWNTO 0); --ADDRESS REG 2
	SIGNAL WB_WR_REG	: STD_LOGIC_VECTOR(4 DOWNTO 0); --WRITE ADDRESS COMING FROM WB STAGE
	SIGNAL WB_RegWrite	: STD_LOGIC; --WRITE SIGNAL ENABLE FROM WB
	
	SIGNAL IM_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0); --immediate generator's output
		
	--PIPE STAGE ID/EX IN
	SIGNAL RD_DATA1: STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA READ 1
	SIGNAL RD_DATA2: STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA READ 2
	SIGNAL IMM_OUT	: STD_LOGIC_VECTOR(31 DOWNTO 0); --IMMEDIATE OUT
	SIGNAL FUNCT		: STD_LOGIC_VECTOR(3 DOWNTO 0); --FUNCTION BITS
	SIGNAL ID_WR_REG	: STD_LOGIC_VECTOR(4 DOWNTO 0); --DECODE STAGE DESTINATION REG ADDRESS
	SIGNAL ID_RD_REG_1 : STD_LOGIC_VECTOR(4 DOWNTO 0); --DECODE STAGE SOURCE REG ADDRESS 1
	SIGNAL ID_RD_REG_2 : STD_LOGIC_VECTOR(4 DOWNTO 0); --DECODE STAGE SOURCE REG ADDRESS 2
	SIGNAL ID_EX_input	:	STD_LOGIC_VECTOR(158 DOWNTO 0); --OVERALL INPUT FOR THE PIPE STAGE
	
--EXECUTION STAGE
	
	--EXECUTION STAGE IN SIGNALS
	SIGNAL ID_EX_output	: 	STD_LOGIC_VECTOR(158 DOWNTO 0); --OVERALL OUTPUT FOR THE PIPE STAGE
	SIGNAL EX_WB		: STD_LOGIC_VECTOR(2 DOWNTO 0); --FROM CU
	SIGNAL EX_M			: STD_LOGIC_VECTOR(2 DOWNTO 0); --FROM CU
	SIGNAL EX_EX		: STD_LOGIC_VECTOR(5 DOWNTO 0); --FROM CU
	SIGNAL EX_I_ADDR	: STD_LOGIC_VECTOR(31 DOWNTO 0); --PC ADDRESS TO EVENTUALLY COMPUTE BRANCH TARGET ADDRESS
	SIGNAL EX_RD_DATA1: STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA READ FROM REG 1
	SIGNAL EX_RD_DATA2: STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA READ FROM REG 2
	SIGNAL EX_IM_OUT	: STD_LOGIC_VECTOR(31 DOWNTO 0); --IMMEDIATE OUT
	SIGNAL EX_FUNCT	: STD_LOGIC_VECTOR(3 DOWNTO 0); --FUNCTION'S BITS
	SIGNAL EX_WR_REG	: STD_LOGIC_VECTOR(4 DOWNTO 0); --DESTINATION REGISTER ADDRESS
	SIGNAL EX_RD_REG_1 : STD_LOGIC_VECTOR(4 DOWNTO 0); --EXECUTE STAGE SOURCE REG ADDRESS 1
	SIGNAL EX_RD_REG_2 : STD_LOGIC_VECTOR(4 DOWNTO 0); --EXECUTE STAGE SOURCE REG ADDRESS 2
	
	--FORWARD UNIT SIGNALS
	SIGNAL MEM_WR_REG : STD_LOGIC_VECTOR(4 DOWNTO 0); --DESTINATION REGISTER ADDRESS FROM MEMORY STAGE
	SIGNAL MUX_FORWARD_A : STD_LOGIC_VECTOR(1 DOWNTO 0); --MUX SELECTION 1
	SIGNAL MUX_FORWARD_B : STD_LOGIC_VECTOR(1 DOWNTO 0); --MUX SELECTION 2
	
	--EXECUTION STAGE SIGNALS
	SIGNAL EX_JMP_ADDR	: STD_LOGIC_VECTOR(31 DOWNTO 0); --OUTPUT OF THE EVENTUAL JUMP ADDRESS
	SIGNAL Z_flag	: STD_LOGIC; --ZERO FLAG (BEQ TAKEN OR NOT)
	SIGNAL ALU_res	: STD_LOGIC_VECTOR(31 DOWNTO 0); --RESULT OF ALU COMPUTATION

	--PIPE STAGE EX/MEM IN
	SIGNAL EX_MEM_input	:	STD_LOGIC_VECTOR(107 DOWNTO 0); --OVERALL INPUT FOR THE PIPE STAGE		--rifare il conto
	
--MEMORY STAGE
	
	--MEMORY STAGE INPUT SIGNALS
	SIGNAL EX_MEM_output	: 	STD_LOGIC_VECTOR(107 DOWNTO 0); --OVERALL OUTPUT FOR THE PIPE STAGE
	SIGNAL MEM_M_branch		: STD_LOGIC; --SIGNAL FOR BRANCH
	SIGNAL MEM_z_flag		: STD_LOGIC; --SIGNAL FOR BRANCH
	SIGNAL MEM_WB			: STD_LOGIC_VECTOR(2 DOWNTO 0); --SIGNAL FROM CU TO WRITE BACK STAGE (4 BITS UNLESS 5 BECAUSE 1 BIT IS USED FOR FORWARDING UNIT FROM MEM STAGE)
	SIGNAL MEM_ALU_Result		: STD_LOGIC_VECTOR(31 DOWNTO 0); --RESULT OF ALU COMPUTATION
	SIGNAL MEM_MemRead		: STD_LOGIC;
	SIGNAL MEM_MemWrite		: STD_LOGIC;
	SIGNAL MEM_WriteData	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	--PIPE STAGE MEM/WB IN
	SIGNAL MEM_WB_input		:	STD_LOGIC_VECTOR(71 DOWNTO 0); --OVERALL INPUT FOR THE PIPE STAGE
	
--WRITE BACK STAGE

	--WRITE BACK STAGE INPUT SIGNALS
	SIGNAL MEM_WB_output	: 	STD_LOGIC_VECTOR(71 DOWNTO 0); --OVERALL OUTPUT FOR THE PIPE STAGE
	SIGNAL MemToReg		: 	STD_LOGIC; --SIGNAL FOR MUX SELECTION
	SIGNAL WB_ReadData	: 	STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA RED FROM MEMORY
	SIGNAL WB_ALU_Result	: 	STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA FROM ALU
	SIGNAL WB_WR_DATA	: 	STD_LOGIC_VECTOR(31 DOWNTO 0); --MUX OUTPUT --PRIMA ERA 32 BIT, MA MI SEMBRA DEBBA ESSERE 64, DA CHIEDERE
	
--HAZARD DETECTION UNIT SIGNALS
	SIGNAL ID_EX_Mem_Read : STD_LOGIC; --ONLY IF THERE'S A LOAD INSTRUCTION, A NOP IS INSERTED
	SIGNAL IF_ID_Write_HD : STD_LOGIC; --SIGNAL TO TURN OFF THE PIPE STAGE ID/EX
	SIGNAL PC_Write_HD : STD_LOGIC; --SIGNAL TO ACTIVATE OR NOT PC
	SIGNAL MUX_CU_HD : STD_LOGIC; --SIGNAL TO SELECT CONTROL UNIT OUTPUT
	
--BRANCH DETECTION UNIT SIGNALS
	SIGNAL D_BRANCH_DET : STD_LOGIC; --SIGNAL TO INSERT A NOP FROM DECODE STAGE
	SIGNAL EX_BRANCH_DET : STD_LOGIC; --SIGNAL TO INSERT A NOP FROM EXECUTION STAGE
	SIGNAL IF_ID_Write_BD : STD_LOGIC; --SIGNAL TO BLOCK PIPE
	SIGNAL PC_Write_BD : STD_LOGIC; --SIGNAL TO ACTIVATE OR NOT PC
	SIGNAL MUX_CU_BD : STD_LOGIC; --SIGNAL TO SELECT CONTROL UNIT OUTPUT
	
	SIGNAL MUX_CU : STD_LOGIC; --OR BETWEEN MUX_CU_BD AND MUX_CU_HD TO SELECT CU OUTPUT
	
	BEGIN
	--Instruction Fetch stage
	seq: sequencer PORT MAP(JUMP_ADDR, PCSrc, PC_Write, clock, reset, I_ADDR);
	PC_address <= I_ADDR;	--I_ADDR is used also to connect the PC to the IF/ID pipe register
	
	--SE ALMENO UNO DEI DUE E' '0', IL RISULTATO E' A ZERO
	PC_Write <= PC_Write_HD AND	PC_Write_BD;
	--IF_ID_Write <= IF_ID_Write_HD AND IF_ID_Write_BD;
	
	IF_ID_input <= I_ADDR & instruction;
	IF_ID_pipe: pipe_register_IF_ID PORT MAP(IF_ID_input, clock, reset, IF_ID_Write_BD, IF_ID_Write_HD, IF_ID_output);
	-- IF_ID_output <= ID_I_ADDR & ID_instruction;

	ID_I_ADDR <= IF_ID_output(63 DOWNTO 32);
	ID_instruction <= IF_ID_output(31 DOWNTO 0);
	
	--Instruction Decode stage
	RD_REG1 <= ID_instruction(19 DOWNTO 15);
	RD_REG2 <= ID_instruction(24 DOWNTO 20);
	OPCODE <= ID_instruction(6 DOWNTO 0);
	FUNCT <= ID_instruction(30) & ID_instruction(14 DOWNTO 12);
	ID_WR_REG <= ID_instruction(11 DOWNTO 7);
	ID_RD_REG_1 <= ID_instruction(19 DOWNTO 15);
	ID_RD_REG_2 <= ID_instruction(24 DOWNTO 20);
	
	JAL_ADDR <= STD_LOGIC_VECTOR(UNSIGNED(ID_I_ADDR) + 4);
	JAL_REGISTER: JAL_REG PORT MAP(JAL_ADDR, clock, reset, WB(2), WR_DATA_JAL);
	
	WITH JAL_SEL SELECT	--connected to the WB(2) coming from the WB stage
		ID_WR_DATA <= WB_WR_DATA WHEN '0',
							WR_DATA_JAL WHEN OTHERS;
	
	RegisterFile: reg_file PORT MAP(RD_REG1, RD_REG2, WB_WR_REG, ID_WR_DATA, WB_RegWrite, clock, reset, RD_DATA1, RD_DATA2);
	ImmGen: immediate_generator PORT MAP(ID_instruction, IM_OUT);
	
	ID_EX_input <= WB & M & EX & ID_I_ADDR & RD_DATA1 & RD_DATA2 & IM_OUT & FUNCT & ID_WR_REG & ID_RD_REG_1 & ID_RD_REG_2;
	ID_EX_pipe: pipe_register_ID_EX PORT MAP(ID_EX_input, clock, reset, '1', ID_EX_output);
	-- ID_EX_output <= EX_WB & EX_M & EX_EX & EX_I_ADDR & EX_RD_DATA1 & EX_RD_DATA2 & EX_IM_OUT & EX_FUNCT & EX_WR_REG & EX_RD_REG_1 & EX_RD_REG_2;
	
	EX_WB <= ID_EX_output(158 DOWNTO 156);
	EX_M <= ID_EX_output(155 DOWNTO 153);
	EX_EX <= ID_EX_output(152 DOWNTO 147);
	EX_I_ADDR <= ID_EX_output(146 DOWNTO 115);
	EX_RD_DATA1 <= ID_EX_output(114 DOWNTO 83);
	EX_RD_DATA2 <= ID_EX_output(82 DOWNTO 51);
	EX_IM_OUT <= ID_EX_output(50 DOWNTO 19);
	EX_FUNCT <= ID_EX_output(18 DOWNTO 15);
	EX_WR_REG <= ID_EX_output(14 DOWNTO 10);
	EX_RD_REG_1 <= ID_EX_output(9 DOWNTO 5);
	EX_RD_REG_2 <= ID_EX_output(4 DOWNTO 0);
	
	--Execution stage
	ex_stage: execution_stage PORT MAP(EX_EX, MUX_FORWARD_A, MUX_FORWARD_B, EX_I_ADDR, EX_RD_DATA1, EX_RD_DATA2, EX_IM_OUT, MEM_ALU_Result, WB_WR_DATA, EX_FUNCT, EX_JMP_ADDR, z_flag, ALU_res);
	
	EX_MEM_input <= EX_WB & EX_M & EX_JMP_ADDR & z_flag & ALU_res & EX_RD_DATA2 & EX_WR_REG; --3+3+32+
	EX_MEM_pipe: pipe_register_EX_MEM PORT MAP(EX_MEM_input, clock, reset, '1', EX_MEM_output);
	--EX_MEM_output <= MEM_WB & MEM_M_branch & MEM_MemRead & MEM_MemWrite & JUMP_ADDR & MEM_z_flag & MEM_ALU_Result & MEM_WriteData & MEM_WR_REG;
	
	MEM_WB <= EX_MEM_output(107 DOWNTO 105);
	MEM_M_branch <= EX_MEM_output(104);
	MemRead <= EX_MEM_output(103);
	MemWrite <= EX_MEM_output(102);
	JUMP_ADDR <= EX_MEM_output(101 DOWNTO 70);
	MEM_z_flag <= EX_MEM_output(69);
	MEM_ALU_Result <= EX_MEM_output(68 DOWNTO 37);
	WriteData <= EX_MEM_output(36 DOWNTO 5);
	MEM_WR_REG <= EX_MEM_output(4 DOWNTO 0);
	
	data_address <= MEM_ALU_Result(31 DOWNTO 0);
	
	--Mem stage
	PCSrc <= MEM_WB(2) OR (MEM_M_branch AND MEM_z_flag);
	
	MEM_WB_input <= MEM_WB & ReadData & MEM_ALU_Result & MEM_WR_REG;
	MEM_WB_pipe: pipe_register_MEM_WB PORT MAP(MEM_WB_input, clock, reset, '1', MEM_WB_output);
	--MEM_WB_output <= JAL_SEL & WB_RegWrite & MemToReg & WB_ReadData & WB_ALU_Result & WB_WR_REG;
	
	JAL_SEL <= MEM_WB_output(71);
	WB_RegWrite <= MEM_WB_output(70);
	MemToReg <= MEM_WB_output(69);
	WB_ReadData <= MEM_WB_output(68 DOWNTO 37);
	WB_ALU_Result <= MEM_WB_output(36 DOWNTO 5);
	WB_WR_REG <= MEM_WB_output(4 DOWNTO 0);
	
	--WB stage
	WITH MemToReg SELECT
	WB_WR_DATA <= WB_ALU_Result when '0',
				  WB_ReadData when OTHERS;
				  
	--FORWARDING unit
	forwarding: forwarding_unit PORT MAP(EX_RD_REG_1, EX_RD_REG_2, MEM_WR_REG, WB_WR_REG, MEM_WB(1), WB_RegWrite, MUX_FORWARD_A, MUX_FORWARD_B);
	
	--HAZARD detection unit
	HDU : hazard_detection_unit PORT MAP(RD_REG1, RD_REG2, EX_WR_REG, EX_M(1), IF_ID_Write_HD, PC_Write_HD, MUX_CU_HD);

	--BRANCH detection unit
	BDU : Branch_Detection PORT MAP(PREMUX_M(2), EX_M(2), PC_Write_BD, IF_ID_Write_BD, MUX_CU_BD);
	
	MUX_CU <= MUX_CU_BD OR MUX_CU_HD;
	
	--Control unit
	CU: control_unit PORT MAP(OPCODE, PREMUX_WB, PREMUX_M, PREMUX_EX);
	WITH MUX_CU SELECT
		 WB <= PREMUX_WB when '0',
			   (OTHERS => '0') when OTHERS;
	WITH MUX_CU SELECT
		 M <= PREMUX_M when '0',
			   (OTHERS => '0') when OTHERS;
	WITH MUX_CU SELECT
		 EX <= PREMUX_EX when '0',
			   (OTHERS => '0') when OTHERS;
END ARCHITECTURE;