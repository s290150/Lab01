Library ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY forwarding_unit IS
	PORT( EX_RS1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			EX_RS2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			MEM_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			WB_RD  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			MEM_SW_BEQ : IN STD_LOGIC; --SE ABBIAMO UNA BEQ O SW NON ABBIAMO REGISTRI DI DESTINAZIONE
			WB_SW_BEQ : IN STD_LOGIC; --SE ABBIAMO UNA BEQ O SW NON ABBIAMO REGISTRI DI DESTINAZIONE
			FORWARD_A : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			FORWARD_B : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEHAVIOUR OF forwarding_unit IS

	SIGNAL forwardA : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL forwardB : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');

BEGIN


	MUX_SELECTION : PROCESS(EX_RS1, EX_RS2, MEM_RD, WB_RD, MEM_SW_BEQ, WB_SW_BEQ)
	BEGIN
		IF ( (MEM_SW_BEQ = '1') AND (WB_SW_BEQ = '1') ) THEN
			IF ( MEM_RD = EX_RS1 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE CICLO PRECEDENTE
				forwardA <= "01";
			ELSIF (  WB_RD = EX_RS1 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE DI DUE CICLI PRIMA
				forwardA <= "10";
			ELSE
				forwardA <= "00";
			END IF;
			IF ( MEM_RD = EX_RS2 ) THEN --DATA DEPENDENCY PER RS2 DA ISTRUZIONE CICLO PRECEDENTE
				forwardB <= "01";
			ELSIF (  WB_RD = EX_RS2 ) THEN --DATA DEPENDENCY PER RS2 DA ISTRUZIONE DI DUE CICLI PRIMA
				forwardB <= "10";
			ELSE
				forwardB <= "00";
			END IF;
		ELSIF ( (MEM_SW_BEQ = '1') AND (WB_SW_BEQ = '0') ) THEN
			IF ( MEM_RD = EX_RS1 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE CICLO PRECEDENTE
				forwardA <= "01";
			ELSE
				forwardA <= "00";
			END IF;
			IF ( MEM_RD = EX_RS2 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE CICLO PRECEDENTE
				forwardB <= "01";
			ELSE
				forwardB <= "00";
			END IF;
		ELSIF ( (MEM_SW_BEQ = '0') AND (WB_SW_BEQ = '1') ) THEN
			IF ( WB_RD = EX_RS1 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE CICLO PRECEDENTE
				forwardA <= "10";
			ELSE
				forwardA <= "00";
			END IF;
			IF ( WB_RD = EX_RS2 ) THEN --DATA DEPENDENCY PER RS1 DA ISTRUZIONE CICLO PRECEDENTE
				forwardB <= "10";
			ELSE
				forwardB <= "00";
			END IF;
		ELSIF ( (MEM_SW_BEQ = '0') AND (WB_SW_BEQ = '0') ) THEN
			forwardA <= "00";
			forwardB <= "00";
		END IF;
	END PROCESS;
	
	
	FORWARD_A <= forwardA;
	FORWARD_B <= forwardB;
	
END ARCHITECTURE;